library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 15;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
  constant RET  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin      

  tmp(0) :=     LDI & "00" & '0' & x"00";
  tmp(1) := 	LDI & "01" & '0' & x"00";
  tmp(2) := 	LDI & "10" & '0' & x"00";
  tmp(3) := 	LDI & "11" & '0' & x"00";
  tmp(4) := 	STA & "00" & '1' & x"20";
  tmp(5) := 	STA & "00" & '1' & x"21";
  tmp(6) := 	STA & "00" & '1' & x"22";
  tmp(7) := 	STA & "00" & '1' & x"23";
  tmp(8) := 	STA & "00" & '1' & x"24";
  tmp(9) := 	STA & "00" & '1' & x"25";
  tmp(10) := 	STA & "00" & '1' & x"00";
  tmp(11) := 	STA & "00" & '1' & x"01";
  tmp(12) := 	STA & "00" & '1' & x"02";
  tmp(13) := 	STA & "00" & '0' & x"00";
  tmp(14) := 	STA & "00" & '0' & x"01";
  tmp(15) := 	STA & "00" & '0' & x"02";
  tmp(16) := 	STA & "00" & '0' & x"03";
  tmp(17) := 	LDI & "00" & '0' & x"09";
  tmp(18) := 	STA & "00" & '0' & x"1E";
  tmp(19) := 	STA & "00" & '0' & x"1F";
  tmp(20) := 	STA & "00" & '0' & x"20";
  tmp(21) := 	STA & "00" & '0' & x"21";
  tmp(22) := 	STA & "00" & '0' & x"22";
  tmp(23) := 	STA & "00" & '0' & x"23";
  tmp(24) := 	LDI & "00" & '0' & x"00";
  tmp(25) := 	STA & "00" & '0' & x"0A";
  tmp(26) := 	LDI & "00" & '0' & x"01";
  tmp(27) := 	STA & "00" & '0' & x"0B";
  tmp(28) := 	LDI & "00" & '0' & x"0A";
  tmp(29) := 	STA & "00" & '0' & x"0C";
  tmp(30) := 	LDI & "00" & '0' & x"01";
  tmp(31) := 	STA & "00" & '0' & x"14";
  tmp(32) := 	LDI & "00" & '0' & x"00";
  tmp(33) := 	STA & "00" & '1' & x"FE";
  tmp(34) := 	STA & "00" & '1' & x"FF";
  tmp(35) := 	STA & "00" & '1' & x"64";
  tmp(36) := 	LDA & "01" & '1' & x"60";
  tmp(37) := 	CEQ & "01" & '0' & x"0A";
  tmp(38) := 	JEQ & "00" & '0' & x"29";
  tmp(39) := 	JSR & "00" & '0' & x"79";
  tmp(40) := 	JSR & "00" & '0' & x"AA";
  tmp(41) := 			LDA & "01" & '1' & x"61";
  tmp(42) := 			CEQ & "01" & '0' & x"0A";
  tmp(43) := 			JEQ & "00" & '0' & x"6D";
  tmp(44) := 			STA & "00" & '1' & x"FE";
  tmp(45) := 				LDI & "00" & '0' & x"01";
  tmp(46) := 				STA & "00" & '1' & x"00";
  tmp(47) := 					LDA & "01" & '1' & x"40";
  tmp(48) := 					STA & "01" & '1' & x"20";
  tmp(49) := 					LDA & "01" & '1' & x"61";
  tmp(50) := 					CEQ & "01" & '0' & x"0A";
  tmp(51) := 					JEQ & "00" & '0' & x"2F";
  tmp(52) := 					STA & "00" & '1' & x"FE";
  tmp(53) := 					STA & "01" & '0' & x"1E";
  tmp(54) := 				LDI & "00" & '0' & x"02";
  tmp(55) := 				STA & "00" & '1' & x"00";
  tmp(56) := 					LDA & "01" & '1' & x"40";
  tmp(57) := 					STA & "01" & '1' & x"21";
  tmp(58) := 					LDA & "01" & '1' & x"61";
  tmp(59) := 					CEQ & "01" & '0' & x"0A";
  tmp(60) := 					JEQ & "00" & '0' & x"38";
  tmp(61) := 					STA & "00" & '1' & x"FE";
  tmp(62) := 					STA & "01" & '0' & x"1F";
  tmp(63) := 				LDI & "00" & '0' & x"04";
  tmp(64) := 				STA & "00" & '1' & x"00";
  tmp(65) := 					LDA & "01" & '1' & x"40";
  tmp(66) := 					STA & "01" & '1' & x"22";
  tmp(67) := 					LDA & "01" & '1' & x"61";
  tmp(68) := 					CEQ & "01" & '0' & x"0A";
  tmp(69) := 					JEQ & "00" & '0' & x"41";
  tmp(70) := 					STA & "00" & '1' & x"FE";
  tmp(71) := 					STA & "01" & '0' & x"20";
  tmp(72) := 				LDI & "00" & '0' & x"08";
  tmp(73) := 				STA & "00" & '1' & x"00";
  tmp(74) := 					LDA & "01" & '1' & x"40";
  tmp(75) := 					STA & "01" & '1' & x"23";
  tmp(76) := 					LDA & "01" & '1' & x"61";
  tmp(77) := 					CEQ & "01" & '0' & x"0A";
  tmp(78) := 					JEQ & "00" & '0' & x"4A";
  tmp(79) := 					STA & "00" & '1' & x"FE";
  tmp(80) := 					STA & "01" & '0' & x"21";
  tmp(81) := 				LDI & "00" & '0' & x"10";
  tmp(82) := 				STA & "00" & '1' & x"00";
  tmp(83) := 					LDA & "01" & '1' & x"40";
  tmp(84) := 					STA & "01" & '1' & x"24";
  tmp(85) := 					LDA & "01" & '1' & x"61";
  tmp(86) := 					CEQ & "01" & '0' & x"0A";
  tmp(87) := 					JEQ & "00" & '0' & x"53";
  tmp(88) := 					STA & "00" & '1' & x"FE";
  tmp(89) := 					STA & "01" & '0' & x"22";
  tmp(90) := 				LDI & "00" & '0' & x"20";
  tmp(91) := 				STA & "00" & '1' & x"00";
  tmp(92) := 					LDA & "01" & '1' & x"40";
  tmp(93) := 					STA & "01" & '1' & x"25";
  tmp(94) := 					LDA & "01" & '1' & x"61";
  tmp(95) := 					CEQ & "01" & '0' & x"0A";
  tmp(96) := 					JEQ & "00" & '0' & x"5C";
  tmp(97) := 					STA & "00" & '1' & x"FE";
  tmp(98) := 					STA & "01" & '0' & x"23";
  tmp(99) := 					LDI & "00" & '0' & x"00";
  tmp(100) := 					LDI & "01" & '0' & x"00";
  tmp(101) := 					STA & "00" & '1' & x"00";
  tmp(102) := 					LDI & "00" & '0' & x"00";
  tmp(103) := 					STA & "00" & '1' & x"20";
  tmp(104) := 					STA & "00" & '1' & x"21";
  tmp(105) := 					STA & "00" & '1' & x"22";
  tmp(106) := 					STA & "00" & '1' & x"23";
  tmp(107) := 					STA & "00" & '1' & x"24";
  tmp(108) := 					STA & "00" & '1' & x"25";
  tmp(109) := 				NOP & "00" & '0' & x"00";
  tmp(110) := JMP  & "00" & '0' & x"24";
  tmp(111) := 	LDI & "10" & '0' & x"00";
  tmp(112) := 	STA & "10" & '0' & x"00";
  tmp(113) := 	STA & "10" & '0' & x"01";
  tmp(114) := 	STA & "10" & '0' & x"02";
  tmp(115) := 	STA & "10" & '0' & x"03";
  tmp(116) := 	STA & "10" & '1' & x"02";
  tmp(117) := 	LDI & "11" & '0' & x"01";
  tmp(118) := 	STA & "11" & '0' & x"14";
  tmp(119) := 	LDI & "11" & '0' & x"00";
  tmp(120) := 	RET & "00" & '0' & x"00";
  tmp(121) := 	STA & "00" & '1' & x"FF";
  tmp(122) := 	LDA & "01" & '0' & x"14";
  tmp(123) := 	CEQ & "01" & '0' & x"0B";
  tmp(124) := 	JEQ & "00" & '0' & x"7E";
  tmp(125) := 	RET & "00" & '0' & x"00";
  tmp(126) := 		SOMA & "10" & '0' & x"0B";
  tmp(127) := 		CEQ & "10" & '0' & x"0C";
  tmp(128) := 		JEQ & "00" & '0' & x"82";
  tmp(129) := 		RET & "00" & '0' & x"00";
  tmp(130) := 			SOMA & "11" & '0' & x"0B";
  tmp(131) := 			CEQ & "11" & '0' & x"0C";
  tmp(132) := 			LDI & "10" & '0' & x"00";
  tmp(133) := 			JEQ & "00" & '0' & x"87";
  tmp(134) := 			RET & "00" & '0' & x"00";
  tmp(135) := 				LDI & "00" & '0' & x"01";
  tmp(136) := 				SOMA & "00" & '0' & x"00";
  tmp(137) := 				LDI & "11" & '0' & x"00";
  tmp(138) := 				CEQ & "00" & '0' & x"0C";
  tmp(139) := 				JEQ & "00" & '0' & x"8E";
  tmp(140) := 				STA & "00" & '0' & x"00";
  tmp(141) := 				RET & "00" & '0' & x"00";
  tmp(142) := 					LDI & "00" & '0' & x"00";
  tmp(143) := 					STA & "00" & '0' & x"00";
  tmp(144) := 					LDI & "00" & '0' & x"01";
  tmp(145) := 					SOMA & "00" & '0' & x"01";
  tmp(146) := 					CEQ & "00" & '0' & x"0C";
  tmp(147) := 					JEQ & "00" & '0' & x"96";
  tmp(148) := 					STA & "00" & '0' & x"01";
  tmp(149) := 					RET & "00" & '0' & x"00";
  tmp(150) := 						LDI & "00" & '0' & x"00";
  tmp(151) := 						STA & "00" & '0' & x"01";
  tmp(152) := 						LDI & "00" & '0' & x"01";
  tmp(153) := 						SOMA & "00" & '0' & x"02";
  tmp(154) := 						CEQ & "00" & '0' & x"0C";
  tmp(155) := 						JEQ & "00" & '0' & x"9E";
  tmp(156) := 						STA & "00" & '0' & x"02";
  tmp(157) := 						RET & "00" & '0' & x"00";
  tmp(158) := 							LDI & "00" & '0' & x"00";
  tmp(159) := 							STA & "00" & '0' & x"02";
  tmp(160) := 							LDI & "00" & '0' & x"01";
  tmp(161) := 							SOMA & "00" & '0' & x"03";
  tmp(162) := 							CEQ & "00" & '0' & x"0C";
  tmp(163) := 							JEQ & "00" & '0' & x"A5";
  tmp(164) := 							RET & "00" & '0' & x"00";
  tmp(165) := 								LDI & "00" & '0' & x"01";
  tmp(166) := 								STA & "00" & '1' & x"02";
  tmp(167) := 								LDI & "00" & '0' & x"00";
  tmp(168) := 								STA & "00" & '0' & x"14";
  tmp(169) := 								RET & "00" & '0' & x"00";
  tmp(170) := 	STA & "10" & '1' & x"20";
  tmp(171) := 	STA & "11" & '1' & x"21";
  tmp(172) := 	LDA & "01" & '0' & x"00";
  tmp(173) := 	STA & "01" & '1' & x"22";
  tmp(174) := 	LDA & "01" & '0' & x"01";
  tmp(175) := 	STA & "01" & '1' & x"23";
  tmp(176) := 	LDA & "01" & '0' & x"02";
  tmp(177) := 	STA & "01" & '1' & x"24";
  tmp(178) := 	LDA & "01" & '0' & x"03";
  tmp(179) := 	STA & "01" & '1' & x"25";
  tmp(180) := 	RET & "00" & '0' & x"00";

        
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;