library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 15;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
  constant RET  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
  constant CLT  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1011";
  constant JLT  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1100";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin      

  tmp(0) :=     LDI & "00" & '0' & x"00";
  tmp(1) := 	LDI & "01" & '0' & x"00";
  tmp(2) := 	LDI & "10" & '0' & x"00";
  tmp(3) := 	LDI & "11" & '0' & x"00";
  tmp(4) := 	STA & "00" & '1' & x"20";
  tmp(5) := 	STA & "00" & '1' & x"21";
  tmp(6) := 	STA & "00" & '1' & x"22";
  tmp(7) := 	STA & "00" & '1' & x"23";
  tmp(8) := 	STA & "00" & '1' & x"24";
  tmp(9) := 	STA & "00" & '1' & x"25";
  tmp(10) := 	STA & "00" & '1' & x"00";
  tmp(11) := 	STA & "00" & '1' & x"01";
  tmp(12) := 	STA & "00" & '1' & x"02";
  tmp(13) := 	STA & "00" & '0' & x"00";
  tmp(14) := 	STA & "00" & '0' & x"01";
  tmp(15) := 	STA & "00" & '0' & x"02";
  tmp(16) := 	STA & "00" & '0' & x"03";
  tmp(17) := 	LDI & "00" & '0' & x"09";
  tmp(18) := 	STA & "00" & '0' & x"1E";
  tmp(19) := 	STA & "00" & '0' & x"1F";
  tmp(20) := 	STA & "00" & '0' & x"20";
  tmp(21) := 	STA & "00" & '0' & x"21";
  tmp(22) := 	STA & "00" & '0' & x"22";
  tmp(23) := 	STA & "00" & '0' & x"23";
  tmp(24) := 	LDI & "00" & '0' & x"00";
  tmp(25) := 	STA & "00" & '0' & x"0A";
  tmp(26) := 	LDI & "00" & '0' & x"01";
  tmp(27) := 	STA & "00" & '0' & x"0B";
  tmp(28) := 	LDI & "00" & '0' & x"0A";
  tmp(29) := 	STA & "00" & '0' & x"0C";
  tmp(30) := 	LDI & "00" & '0' & x"06";
  tmp(31) := 	STA & "00" & '0' & x"0D";
  tmp(32) := 	LDI & "00" & '0' & x"04";
  tmp(33) := 	STA & "00" & '0' & x"0E";
  tmp(34) := 	LDI & "00" & '0' & x"02";
  tmp(35) := 	STA & "00" & '0' & x"0F";
  tmp(36) := 	LDI & "00" & '0' & x"01";
  tmp(37) := 	STA & "00" & '0' & x"14";
  tmp(38) := 	LDI & "00" & '0' & x"01";
  tmp(39) := 	STA & "00" & '0' & x"15";
  tmp(40) := 	LDI & "00" & '0' & x"00";
  tmp(41) := 	STA & "00" & '0' & x"16";
  tmp(42) := 	LDI & "00" & '0' & x"00";
  tmp(43) := 	STA & "00" & '1' & x"FE";
  tmp(44) := 	STA & "00" & '1' & x"FC";
  tmp(45) := 	STA & "00" & '1' & x"FD";
  tmp(46) := 	LDA & "01" & '1' & x"65";
  tmp(47) := 	CEQ & "01" & '0' & x"0A";
  tmp(48) := 	JSR & "00" & '1' & x"4B";
  tmp(49) := 	JEQ & "00" & '0' & x"37";
  tmp(50) := 	JSR & "00" & '0' & x"FC";
  tmp(51) := 	LDA & "01" & '1' & x"64";
  tmp(52) := 	CEQ & "01" & '0' & x"0A";
  tmp(53) := 	JEQ & "00" & '0' & x"37";
  tmp(54) := 	JSR & "00" & '0' & x"EA";
  tmp(55) := 			LDA & "01" & '1' & x"61";
  tmp(56) := 			CEQ & "01" & '0' & x"0A";
  tmp(57) := 			JEQ & "00" & '0' & x"3B";
  tmp(58) := 			STA & "00" & '1' & x"FE";
  tmp(59) := 				STA & "00" & '1' & x"FE";
  tmp(60) := 				LDA & "01" & '1' & x"60";
  tmp(61) := 				CEQ & "01" & '0' & x"0A";
  tmp(62) := 				JEQ & "00" & '0' & x"40";
  tmp(63) := 				JSR & "00" & '0' & x"43";
  tmp(64) := 					NOP & "00" & '0' & x"00";
  tmp(65) := JMP  & "00" & '0' & x"2E";
  tmp(66) := STA  & "00" & '0' & x"00";
  tmp(67) := 	LDI & "00" & '0' & x"00";
  tmp(68) := 	STA & "00" & '1' & x"20";
  tmp(69) := 	STA & "00" & '1' & x"21";
  tmp(70) := 	STA & "00" & '1' & x"22";
  tmp(71) := 	STA & "00" & '1' & x"23";
  tmp(72) := 	STA & "00" & '1' & x"24";
  tmp(73) := 	STA & "00" & '1' & x"25";
  tmp(74) := STA  & "00" & '0' & x"00";
  tmp(75) := 		STA & "00" & '1' & x"FF";
  tmp(76) := 		LDI & "00" & '0' & x"01";
  tmp(77) := 		STA & "00" & '1' & x"02";
  tmp(78) := 			LDA & "00" & '1' & x"40";
  tmp(79) := 			LDA & "01" & '0' & x"15";
  tmp(80) := 			CEQ & "01" & '0' & x"0A";
  tmp(81) := 			JEQ & "00" & '0' & x"5E";
  tmp(82) := 			LDI & "01" & '0' & x"02";
  tmp(83) := 			CLT & "01" & '1' & x"40";
  tmp(84) := 			JLT & "00" & '0' & x"56";
  tmp(85) := 			JMP & "00" & '0' & x"57";
  tmp(86) := 				LDI & "00" & '0' & x"02";
  tmp(87) := 				STA & "00" & '1' & x"25";
  tmp(88) := 				LDA & "01" & '1' & x"60";
  tmp(89) := 				CEQ & "01" & '0' & x"0A";
  tmp(90) := 				JEQ & "00" & '0' & x"4E";
  tmp(91) := 				STA & "00" & '1' & x"FF";
  tmp(92) := 				STA & "00" & '0' & x"03";
  tmp(93) := 				JMP & "00" & '0' & x"6A";
  tmp(94) := 				LDI & "01" & '0' & x"01";
  tmp(95) := 				CLT & "01" & '1' & x"40";
  tmp(96) := 				JLT & "00" & '0' & x"62";
  tmp(97) := 				JMP & "00" & '0' & x"63";
  tmp(98) := 					LDI & "00" & '0' & x"01";
  tmp(99) := 					STA & "00" & '1' & x"25";
  tmp(100) := 					LDA & "01" & '1' & x"60";
  tmp(101) := 					CEQ & "01" & '0' & x"0A";
  tmp(102) := 					JEQ & "00" & '0' & x"4E";
  tmp(103) := 					STA & "00" & '1' & x"FF";
  tmp(104) := 					STA & "00" & '0' & x"03";
  tmp(105) := STA  & "00" & '0' & x"00";
  tmp(106) := 		STA & "00" & '1' & x"FF";
  tmp(107) := 		LDI & "00" & '0' & x"01";
  tmp(108) := 		STA & "00" & '1' & x"01";
  tmp(109) := 			LDA & "00" & '1' & x"40";
  tmp(110) := 			LDA & "01" & '0' & x"15";
  tmp(111) := 			CEQ & "01" & '0' & x"0A";
  tmp(112) := 			JEQ & "00" & '0' & x"8C";
  tmp(113) := 			LDI & "01" & '0' & x"02";
  tmp(114) := 			CEQ & "01" & '0' & x"03";
  tmp(115) := 			JEQ & "00" & '0' & x"80";
  tmp(116) := 			LDI & "01" & '0' & x"0A";
  tmp(117) := 			CLT & "01" & '1' & x"40";
  tmp(118) := 			JLT & "00" & '0' & x"78";
  tmp(119) := 			JMP & "00" & '0' & x"79";
  tmp(120) := 				LDI & "00" & '0' & x"09";
  tmp(121) := 				STA & "00" & '1' & x"24";
  tmp(122) := 				LDA & "01" & '1' & x"60";
  tmp(123) := 				CEQ & "01" & '0' & x"0A";
  tmp(124) := 				JEQ & "00" & '0' & x"6D";
  tmp(125) := 				STA & "00" & '1' & x"FF";
  tmp(126) := 				STA & "00" & '0' & x"02";
  tmp(127) := 				JMP & "00" & '0' & x"A7";
  tmp(128) := 				LDI & "01" & '0' & x"03";
  tmp(129) := 				CLT & "01" & '1' & x"40";
  tmp(130) := 				JLT & "00" & '0' & x"84";
  tmp(131) := 				JMP & "00" & '0' & x"85";
  tmp(132) := 					LDI & "00" & '0' & x"03";
  tmp(133) := 					STA & "00" & '1' & x"24";
  tmp(134) := 					LDA & "01" & '1' & x"60";
  tmp(135) := 					CEQ & "01" & '0' & x"0A";
  tmp(136) := 					JEQ & "00" & '0' & x"6D";
  tmp(137) := 					STA & "00" & '1' & x"FF";
  tmp(138) := 					STA & "00" & '0' & x"02";
  tmp(139) := 					JMP & "00" & '0' & x"A7";
  tmp(140) := 				LDI & "01" & '0' & x"01";
  tmp(141) := 				CEQ & "01" & '0' & x"03";
  tmp(142) := 				JEQ & "00" & '0' & x"9B";
  tmp(143) := 				LDI & "01" & '0' & x"0A";
  tmp(144) := 				CLT & "01" & '1' & x"40";
  tmp(145) := 				JLT & "00" & '0' & x"93";
  tmp(146) := 				JMP & "00" & '0' & x"94";
  tmp(147) := 					LDI & "00" & '0' & x"09";
  tmp(148) := 					STA & "00" & '1' & x"24";
  tmp(149) := 					LDA & "01" & '1' & x"60";
  tmp(150) := 					CEQ & "01" & '0' & x"0A";
  tmp(151) := 					JEQ & "00" & '0' & x"6D";
  tmp(152) := 					STA & "00" & '1' & x"FF";
  tmp(153) := 					STA & "00" & '0' & x"02";
  tmp(154) := 					JMP & "00" & '0' & x"A7";
  tmp(155) := 					LDI & "01" & '0' & x"02";
  tmp(156) := 					CLT & "01" & '1' & x"40";
  tmp(157) := 					JLT & "00" & '0' & x"9F";
  tmp(158) := 					JMP & "00" & '0' & x"A0";
  tmp(159) := 						LDI & "00" & '0' & x"01";
  tmp(160) := 						STA & "00" & '1' & x"24";
  tmp(161) := 						LDA & "01" & '1' & x"60";
  tmp(162) := 						CEQ & "01" & '0' & x"0A";
  tmp(163) := 						JEQ & "00" & '0' & x"6D";
  tmp(164) := 						STA & "00" & '1' & x"FF";
  tmp(165) := 						STA & "00" & '0' & x"02";
  tmp(166) := STA  & "00" & '0' & x"00";
  tmp(167) := 		STA & "00" & '1' & x"FF";
  tmp(168) := 		LDI & "00" & '0' & x"80";
  tmp(169) := 		STA & "00" & '1' & x"00";
  tmp(170) := 			LDA & "00" & '1' & x"40";
  tmp(171) := 			LDI & "01" & '0' & x"06";
  tmp(172) := 			CLT & "01" & '1' & x"40";
  tmp(173) := 			JLT & "00" & '0' & x"AF";
  tmp(174) := 			JMP & "00" & '0' & x"B0";
  tmp(175) := 				LDI & "00" & '0' & x"05";
  tmp(176) := 				STA & "00" & '1' & x"23";
  tmp(177) := 				LDA & "01" & '1' & x"60";
  tmp(178) := 				CEQ & "01" & '0' & x"0A";
  tmp(179) := 				JEQ & "00" & '0' & x"AA";
  tmp(180) := 				STA & "00" & '1' & x"FF";
  tmp(181) := 				STA & "00" & '0' & x"01";
  tmp(182) := STA  & "00" & '0' & x"00";
  tmp(183) := 		STA & "00" & '1' & x"FF";
  tmp(184) := 		LDI & "00" & '0' & x"C0";
  tmp(185) := 		STA & "00" & '1' & x"00";
  tmp(186) := 			LDA & "00" & '1' & x"40";
  tmp(187) := 			LDI & "01" & '0' & x"0A";
  tmp(188) := 			CLT & "01" & '1' & x"40";
  tmp(189) := 			JLT & "00" & '0' & x"BF";
  tmp(190) := 			JMP & "00" & '0' & x"C0";
  tmp(191) := 				LDI & "00" & '0' & x"09";
  tmp(192) := 				STA & "00" & '1' & x"22";
  tmp(193) := 				LDA & "01" & '1' & x"60";
  tmp(194) := 				CEQ & "01" & '0' & x"0A";
  tmp(195) := 				JEQ & "00" & '0' & x"BA";
  tmp(196) := 				STA & "00" & '1' & x"FF";
  tmp(197) := 				STA & "00" & '0' & x"00";
  tmp(198) := STA  & "00" & '0' & x"00";
  tmp(199) := 		STA & "00" & '1' & x"FF";
  tmp(200) := 		LDI & "00" & '0' & x"E0";
  tmp(201) := 		STA & "00" & '1' & x"00";
  tmp(202) := 			LDA & "11" & '1' & x"40";
  tmp(203) := 			LDI & "01" & '0' & x"06";
  tmp(204) := 			CLT & "01" & '1' & x"40";
  tmp(205) := 			JLT & "00" & '0' & x"CF";
  tmp(206) := 			JMP & "00" & '0' & x"D0";
  tmp(207) := 				LDI & "11" & '0' & x"05";
  tmp(208) := 				STA & "11" & '1' & x"21";
  tmp(209) := 				LDA & "01" & '1' & x"60";
  tmp(210) := 				CEQ & "01" & '0' & x"0A";
  tmp(211) := 				JEQ & "00" & '0' & x"CA";
  tmp(212) := 				STA & "00" & '1' & x"FF";
  tmp(213) := STA  & "00" & '0' & x"00";
  tmp(214) := 		STA & "00" & '1' & x"FF";
  tmp(215) := 		LDI & "00" & '0' & x"F0";
  tmp(216) := 		STA & "00" & '1' & x"00";
  tmp(217) := 			LDA & "10" & '1' & x"40";
  tmp(218) := 			LDI & "01" & '0' & x"0A";
  tmp(219) := 			CLT & "01" & '1' & x"40";
  tmp(220) := 			JLT & "00" & '0' & x"DE";
  tmp(221) := 			JMP & "00" & '0' & x"DF";
  tmp(222) := 				LDI & "10" & '0' & x"09";
  tmp(223) := 				STA & "10" & '1' & x"20";
  tmp(224) := 				LDA & "01" & '1' & x"60";
  tmp(225) := 				CEQ & "01" & '0' & x"0A";
  tmp(226) := 				JEQ & "00" & '0' & x"D9";
  tmp(227) := 				STA & "00" & '1' & x"FF";
  tmp(228) := 				LDI & "00" & '0' & x"00";
  tmp(229) := 				LDI & "01" & '0' & x"00";
  tmp(230) := 				STA & "00" & '1' & x"00";
  tmp(231) := 				STA & "00" & '1' & x"01";
  tmp(232) := 				STA & "00" & '1' & x"02";
  tmp(233) := 				RET & "00" & '0' & x"00";
  tmp(234) := 	STA & "00" & '1' & x"FD";
  tmp(235) := 	LDI & "10" & '0' & x"00";
  tmp(236) := 	STA & "10" & '0' & x"00";
  tmp(237) := 	STA & "10" & '0' & x"01";
  tmp(238) := 	STA & "10" & '0' & x"02";
  tmp(239) := 	STA & "10" & '0' & x"03";
  tmp(240) := 	STA & "10" & '1' & x"20";
  tmp(241) := 	STA & "10" & '1' & x"21";
  tmp(242) := 	STA & "10" & '1' & x"22";
  tmp(243) := 	STA & "10" & '1' & x"23";
  tmp(244) := 	STA & "10" & '1' & x"24";
  tmp(245) := 	STA & "10" & '1' & x"25";
  tmp(246) := 	STA & "10" & '1' & x"01";
  tmp(247) := 	STA & "10" & '1' & x"02";
  tmp(248) := 	LDI & "11" & '0' & x"01";
  tmp(249) := 	STA & "11" & '0' & x"14";
  tmp(250) := 	LDI & "11" & '0' & x"00";
  tmp(251) := 	RET & "00" & '0' & x"00";
  tmp(252) := 	STA & "00" & '1' & x"FC";
  tmp(253) := 	LDA & "01" & '0' & x"14";
  tmp(254) := 	CEQ & "01" & '0' & x"0B";
  tmp(255) := 	JEQ & "00" & '1' & x"01";
  tmp(256) := 	RET & "00" & '0' & x"00";
  tmp(257) := 		SOMA & "10" & '0' & x"0B";
  tmp(258) := 		CEQ & "10" & '0' & x"0C";
  tmp(259) := 		JEQ & "00" & '1' & x"05";
  tmp(260) := 		RET & "00" & '0' & x"00";
  tmp(261) := 			SOMA & "11" & '0' & x"0B";
  tmp(262) := 			CEQ & "11" & '0' & x"0D";
  tmp(263) := 			LDI & "10" & '0' & x"00";
  tmp(264) := 			JEQ & "00" & '1' & x"0A";
  tmp(265) := 			RET & "00" & '0' & x"00";
  tmp(266) := 				LDI & "00" & '0' & x"01";
  tmp(267) := 				SOMA & "00" & '0' & x"00";
  tmp(268) := 				LDI & "11" & '0' & x"00";
  tmp(269) := 				CEQ & "00" & '0' & x"0C";
  tmp(270) := 				JEQ & "00" & '1' & x"11";
  tmp(271) := 				STA & "00" & '0' & x"00";
  tmp(272) := 				RET & "00" & '0' & x"00";
  tmp(273) := 					LDI & "00" & '0' & x"00";
  tmp(274) := 					STA & "00" & '0' & x"00";
  tmp(275) := 					LDI & "00" & '0' & x"01";
  tmp(276) := 					SOMA & "00" & '0' & x"01";
  tmp(277) := 					CEQ & "00" & '0' & x"0D";
  tmp(278) := 					JEQ & "00" & '1' & x"19";
  tmp(279) := 					STA & "00" & '0' & x"01";
  tmp(280) := 					RET & "00" & '0' & x"00";
  tmp(281) := 						LDI & "00" & '0' & x"00";
  tmp(282) := 						STA & "00" & '0' & x"01";
  tmp(283) := 						LDI & "00" & '0' & x"01";
  tmp(284) := 						SOMA & "00" & '0' & x"02";
  tmp(285) := 						CEQ & "00" & '0' & x"0C";
  tmp(286) := 						JEQ & "00" & '1' & x"21";
  tmp(287) := 						STA & "00" & '0' & x"02";
  tmp(288) := 						JMP & "00" & '1' & x"26";
  tmp(289) := 							LDI & "00" & '0' & x"00";
  tmp(290) := 							STA & "00" & '0' & x"02";
  tmp(291) := 							LDI & "00" & '0' & x"01";
  tmp(292) := 							SOMA & "00" & '0' & x"03";
  tmp(293) := 							STA & "00" & '0' & x"03";
  tmp(294) := 			LDA & "00" & '0' & x"15";
  tmp(295) := 			CEQ & "00" & '0' & x"0A";
  tmp(296) := 			JEQ & "00" & '1' & x"35";
  tmp(297) := 			LDA & "00" & '0' & x"02";
  tmp(298) := 			CEQ & "00" & '0' & x"0E";
  tmp(299) := 			JEQ & "00" & '1' & x"2D";
  tmp(300) := 			RET & "00" & '0' & x"00";
  tmp(301) := 					LDA & "00" & '0' & x"03";
  tmp(302) := 					CEQ & "00" & '0' & x"0F";
  tmp(303) := 					JEQ & "00" & '1' & x"31";
  tmp(304) := 					RET & "00" & '0' & x"00";
  tmp(305) := 							LDI & "00" & '0' & x"00";
  tmp(306) := 							STA & "00" & '0' & x"02";
  tmp(307) := 							STA & "00" & '0' & x"03";
  tmp(308) := 							RET & "00" & '0' & x"00";
  tmp(309) := 				LDA & "00" & '0' & x"02";
  tmp(310) := 				CEQ & "00" & '0' & x"0F";
  tmp(311) := 				JEQ & "00" & '1' & x"39";
  tmp(312) := 				RET & "00" & '0' & x"00";
  tmp(313) := 						LDA & "00" & '0' & x"03";
  tmp(314) := 						CEQ & "00" & '0' & x"0B";
  tmp(315) := 						JEQ & "00" & '1' & x"3D";
  tmp(316) := 						RET & "00" & '0' & x"00";
  tmp(317) := 								LDI & "00" & '0' & x"00";
  tmp(318) := 								STA & "00" & '0' & x"02";
  tmp(319) := 								STA & "00" & '0' & x"03";
  tmp(320) := 								LDA & "00" & '0' & x"16";
  tmp(321) := 								CEQ & "00" & '0' & x"0A";
  tmp(322) := 								JEQ & "00" & '1' & x"47";
  tmp(323) := 								LDI & "00" & '0' & x"00";
  tmp(324) := 								STA & "00" & '0' & x"16";
  tmp(325) := 								STA & "00" & '1' & x"02";
  tmp(326) := 								RET & "00" & '0' & x"00";
  tmp(327) := 										LDI & "00" & '0' & x"01";
  tmp(328) := 										STA & "00" & '0' & x"16";
  tmp(329) := 										STA & "00" & '1' & x"02";
  tmp(330) := 										RET & "00" & '0' & x"00";
  tmp(331) := 	STA & "10" & '1' & x"20";
  tmp(332) := 	STA & "11" & '1' & x"21";
  tmp(333) := 	LDA & "01" & '0' & x"00";
  tmp(334) := 	STA & "01" & '1' & x"22";
  tmp(335) := 	LDA & "01" & '0' & x"01";
  tmp(336) := 	STA & "01" & '1' & x"23";
  tmp(337) := 	LDA & "01" & '0' & x"02";
  tmp(338) := 	STA & "01" & '1' & x"24";
  tmp(339) := 	LDA & "01" & '0' & x"03";
  tmp(340) := 	STA & "01" & '1' & x"25";
  tmp(341) := 	RET & "00" & '0' & x"00";
        
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;