library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 15;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
  constant RET  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin      

  tmp(0) :=     LDI & "00" & '0' & x"00";
tmp(1) := 	LDI & "01" & '0' & x"00";
tmp(2) := 	LDI & "10" & '0' & x"00";
tmp(3) := 	LDI & "11" & '0' & x"00";
tmp(4) := 	STA & "00" & '1' & x"20";
tmp(5) := 	STA & "00" & '1' & x"21";
tmp(6) := 	STA & "00" & '1' & x"22";
tmp(7) := 	STA & "00" & '1' & x"23";
tmp(8) := 	STA & "00" & '1' & x"24";
tmp(9) := 	STA & "00" & '1' & x"25";
tmp(10) := 	STA & "00" & '1' & x"00";
tmp(11) := 	STA & "00" & '1' & x"01";
tmp(12) := 	STA & "00" & '1' & x"02";
tmp(13) := 	STA & "00" & '0' & x"00";
tmp(14) := 	STA & "00" & '0' & x"01";
tmp(15) := 	STA & "00" & '0' & x"02";
tmp(16) := 	STA & "00" & '0' & x"03";
tmp(17) := 	LDI & "00" & '0' & x"09";
tmp(18) := 	STA & "00" & '0' & x"1E";
tmp(19) := 	STA & "00" & '0' & x"1F";
tmp(20) := 	STA & "00" & '0' & x"20";
tmp(21) := 	STA & "00" & '0' & x"21";
tmp(22) := 	STA & "00" & '0' & x"22";
tmp(23) := 	STA & "00" & '0' & x"23";
tmp(24) := 	LDI & "00" & '0' & x"00";
tmp(25) := 	STA & "00" & '0' & x"0A";
tmp(26) := 	LDI & "00" & '0' & x"01";
tmp(27) := 	STA & "00" & '0' & x"0B";
tmp(28) := 	LDI & "00" & '0' & x"0A";
tmp(29) := 	STA & "00" & '0' & x"0C";
tmp(30) := 	LDI & "00" & '0' & x"06";
tmp(31) := 	STA & "00" & '0' & x"0D";
tmp(32) := 	LDI & "00" & '0' & x"04";
tmp(33) := 	STA & "00" & '0' & x"0E";
tmp(34) := 	LDI & "00" & '0' & x"02";
tmp(35) := 	STA & "00" & '0' & x"0F";
tmp(36) := 	LDI & "00" & '0' & x"01";
tmp(37) := 	STA & "00" & '0' & x"14";
tmp(38) := 	LDI & "00" & '0' & x"00";
tmp(39) := 	STA & "00" & '0' & x"15";
tmp(40) := 	LDI & "00" & '0' & x"00";
tmp(41) := 	STA & "00" & '0' & x"16";
tmp(42) := 	LDI & "00" & '0' & x"00";
tmp(43) := 	STA & "00" & '1' & x"FE";
tmp(44) := 	STA & "00" & '1' & x"FC";
tmp(45) := 	STA & "00" & '1' & x"FD";
tmp(46) := 	LDA & "01" & '1' & x"65";
tmp(47) := 	CEQ & "01" & '0' & x"0A";
tmp(48) := 	JSR & "00" & '0' & x"DF";
tmp(49) := 	JEQ & "00" & '0' & x"38";
tmp(50) := 	JSR & "00" & '0' & x"EA";
tmp(51) := 	JSR & "00" & '0' & x"90";
tmp(52) := 	LDA & "01" & '1' & x"64";
tmp(53) := 	CEQ & "01" & '0' & x"0A";
tmp(54) := 	JEQ & "00" & '0' & x"38";
tmp(55) := 	JSR & "00" & '0' & x"7E";
tmp(56) := 			LDA & "01" & '1' & x"61";
tmp(57) := 			CEQ & "01" & '0' & x"0A";
tmp(58) := 			JEQ & "00" & '0' & x"7C";
tmp(59) := 			STA & "00" & '1' & x"FE";
tmp(60) := 				LDI & "00" & '0' & x"01";
tmp(61) := 				STA & "00" & '1' & x"00";
tmp(62) := 					LDA & "00" & '1' & x"40";
tmp(63) := 					STA & "00" & '1' & x"20";
tmp(64) := 					LDA & "01" & '1' & x"61";
tmp(65) := 					CEQ & "01" & '0' & x"0A";
tmp(66) := 					JEQ & "00" & '0' & x"3E";
tmp(67) := 					STA & "00" & '1' & x"FE";
tmp(68) := 					STA & "00" & '0' & x"1E";
tmp(69) := 				LDI & "00" & '0' & x"02";
tmp(70) := 				STA & "00" & '1' & x"00";
tmp(71) := 					LDA & "00" & '1' & x"40";
tmp(72) := 					STA & "00" & '1' & x"21";
tmp(73) := 					LDA & "01" & '1' & x"61";
tmp(74) := 					CEQ & "01" & '0' & x"0A";
tmp(75) := 					JEQ & "00" & '0' & x"47";
tmp(76) := 					STA & "00" & '1' & x"FE";
tmp(77) := 					STA & "00" & '0' & x"1F";
tmp(78) := 				LDI & "00" & '0' & x"04";
tmp(79) := 				STA & "00" & '1' & x"00";
tmp(80) := 					LDA & "00" & '1' & x"40";
tmp(81) := 					STA & "00" & '1' & x"22";
tmp(82) := 					LDA & "01" & '1' & x"61";
tmp(83) := 					CEQ & "01" & '0' & x"0A";
tmp(84) := 					JEQ & "00" & '0' & x"50";
tmp(85) := 					STA & "00" & '1' & x"FE";
tmp(86) := 					STA & "00" & '0' & x"20";
tmp(87) := 				LDI & "00" & '0' & x"08";
tmp(88) := 				STA & "00" & '1' & x"00";
tmp(89) := 					LDA & "00" & '1' & x"40";
tmp(90) := 					STA & "00" & '1' & x"23";
tmp(91) := 					LDA & "01" & '1' & x"61";
tmp(92) := 					CEQ & "01" & '0' & x"0A";
tmp(93) := 					JEQ & "00" & '0' & x"59";
tmp(94) := 					STA & "00" & '1' & x"FE";
tmp(95) := 					STA & "00" & '0' & x"21";
tmp(96) := 				LDI & "00" & '0' & x"10";
tmp(97) := 				STA & "00" & '1' & x"00";
tmp(98) := 					LDA & "00" & '1' & x"40";
tmp(99) := 					STA & "00" & '1' & x"24";
tmp(100) := 					LDA & "01" & '1' & x"61";
tmp(101) := 					CEQ & "01" & '0' & x"0A";
tmp(102) := 					JEQ & "00" & '0' & x"62";
tmp(103) := 					STA & "00" & '1' & x"FE";
tmp(104) := 					STA & "00" & '0' & x"22";
tmp(105) := 				LDI & "00" & '0' & x"20";
tmp(106) := 				STA & "00" & '1' & x"00";
tmp(107) := 					LDA & "00" & '1' & x"40";
tmp(108) := 					STA & "00" & '1' & x"25";
tmp(109) := 					LDA & "01" & '1' & x"61";
tmp(110) := 					CEQ & "01" & '0' & x"0A";
tmp(111) := 					JEQ & "00" & '0' & x"6B";
tmp(112) := 					STA & "00" & '1' & x"FE";
tmp(113) := 					STA & "00" & '0' & x"23";
tmp(114) := 					LDI & "00" & '0' & x"00";
tmp(115) := 					LDI & "01" & '0' & x"00";
tmp(116) := 					STA & "00" & '1' & x"00";
tmp(117) := 					LDI & "00" & '0' & x"00";
tmp(118) := 					STA & "00" & '1' & x"20";
tmp(119) := 					STA & "00" & '1' & x"21";
tmp(120) := 					STA & "00" & '1' & x"22";
tmp(121) := 					STA & "00" & '1' & x"23";
tmp(122) := 					STA & "00" & '1' & x"24";
tmp(123) := 					STA & "00" & '1' & x"25";
tmp(124) := 				NOP & "00" & '0' & x"00";
tmp(125) := JMP  & "00" & '0' & x"2E";
tmp(126) := 	STA & "00" & '1' & x"FD";
tmp(127) := 	LDI & "10" & '0' & x"00";
tmp(128) := 	STA & "10" & '0' & x"00";
tmp(129) := 	STA & "10" & '0' & x"01";
tmp(130) := 	STA & "10" & '0' & x"02";
tmp(131) := 	STA & "10" & '0' & x"03";
tmp(132) := 	STA & "10" & '1' & x"20";
tmp(133) := 	STA & "10" & '1' & x"21";
tmp(134) := 	STA & "10" & '1' & x"22";
tmp(135) := 	STA & "10" & '1' & x"23";
tmp(136) := 	STA & "10" & '1' & x"24";
tmp(137) := 	STA & "10" & '1' & x"25";
tmp(138) := 	STA & "10" & '1' & x"01";
tmp(139) := 	STA & "10" & '1' & x"02";
tmp(140) := 	LDI & "11" & '0' & x"01";
tmp(141) := 	STA & "11" & '0' & x"14";
tmp(142) := 	LDI & "11" & '0' & x"00";
tmp(143) := 	RET & "00" & '0' & x"00";
tmp(144) := 	STA & "00" & '1' & x"FC";
tmp(145) := 	LDA & "01" & '0' & x"14";
tmp(146) := 	CEQ & "01" & '0' & x"0B";
tmp(147) := 	JEQ & "00" & '0' & x"95";
tmp(148) := 	RET & "00" & '0' & x"00";
tmp(149) := 		SOMA & "10" & '0' & x"0B";
tmp(150) := 		CEQ & "10" & '0' & x"0C";
tmp(151) := 		JEQ & "00" & '0' & x"99";
tmp(152) := 		RET & "00" & '0' & x"00";
tmp(153) := 			SOMA & "11" & '0' & x"0B";
tmp(154) := 			CEQ & "11" & '0' & x"0D";
tmp(155) := 			LDI & "10" & '0' & x"00";
tmp(156) := 			JEQ & "00" & '0' & x"9E";
tmp(157) := 			RET & "00" & '0' & x"00";
tmp(158) := 				LDI & "00" & '0' & x"01";
tmp(159) := 				SOMA & "00" & '0' & x"00";
tmp(160) := 				LDI & "11" & '0' & x"00";
tmp(161) := 				CEQ & "00" & '0' & x"0C";
tmp(162) := 				JEQ & "00" & '0' & x"A5";
tmp(163) := 				STA & "00" & '0' & x"00";
tmp(164) := 				RET & "00" & '0' & x"00";
tmp(165) := 					LDI & "00" & '0' & x"00";
tmp(166) := 					STA & "00" & '0' & x"00";
tmp(167) := 					LDI & "00" & '0' & x"01";
tmp(168) := 					SOMA & "00" & '0' & x"01";
tmp(169) := 					CEQ & "00" & '0' & x"0D";
tmp(170) := 					JEQ & "00" & '0' & x"AD";
tmp(171) := 					STA & "00" & '0' & x"01";
tmp(172) := 					RET & "00" & '0' & x"00";
tmp(173) := 						LDI & "00" & '0' & x"00";
tmp(174) := 						STA & "00" & '0' & x"01";
tmp(175) := 						LDI & "00" & '0' & x"01";
tmp(176) := 						SOMA & "00" & '0' & x"02";
tmp(177) := 						CEQ & "00" & '0' & x"0C";
tmp(178) := 						JEQ & "00" & '0' & x"B5";
tmp(179) := 						STA & "00" & '0' & x"02";
tmp(180) := 						JMP & "00" & '0' & x"BA";
tmp(181) := 							LDI & "00" & '0' & x"00";
tmp(182) := 							STA & "00" & '0' & x"02";
tmp(183) := 							LDI & "00" & '0' & x"01";
tmp(184) := 							SOMA & "00" & '0' & x"03";
tmp(185) := 							STA & "00" & '0' & x"03";
tmp(186) := 			LDA & "00" & '0' & x"15";
tmp(187) := 			CEQ & "00" & '0' & x"0A";
tmp(188) := 			JEQ & "00" & '0' & x"C9";
tmp(189) := 			LDA & "00" & '0' & x"02";
tmp(190) := 			CEQ & "00" & '0' & x"0E";
tmp(191) := 			JEQ & "00" & '0' & x"C1";
tmp(192) := 			RET & "00" & '0' & x"00";
tmp(193) := 					LDA & "00" & '0' & x"03";
tmp(194) := 					CEQ & "00" & '0' & x"0F";
tmp(195) := 					JEQ & "00" & '0' & x"C5";
tmp(196) := 					RET & "00" & '0' & x"00";
tmp(197) := 							LDI & "00" & '0' & x"00";
tmp(198) := 							STA & "00" & '0' & x"02";
tmp(199) := 							STA & "00" & '0' & x"03";
tmp(200) := 							RET & "00" & '0' & x"00";
tmp(201) := 				LDA & "00" & '0' & x"02";
tmp(202) := 				CEQ & "00" & '0' & x"0F";
tmp(203) := 				JEQ & "00" & '0' & x"CD";
tmp(204) := 				RET & "00" & '0' & x"00";
tmp(205) := 						LDA & "00" & '0' & x"03";
tmp(206) := 						CEQ & "00" & '0' & x"0B";
tmp(207) := 						JEQ & "00" & '0' & x"D1";
tmp(208) := 						RET & "00" & '0' & x"00";
tmp(209) := 								LDI & "00" & '0' & x"00";
tmp(210) := 								STA & "00" & '0' & x"02";
tmp(211) := 								STA & "00" & '0' & x"03";
tmp(212) := 								LDA & "00" & '0' & x"16";
tmp(213) := 								CEQ & "00" & '0' & x"0A";
tmp(214) := 								JEQ & "00" & '0' & x"DB";
tmp(215) := 								LDI & "00" & '0' & x"00";
tmp(216) := 								STA & "00" & '0' & x"16";
tmp(217) := 								STA & "00" & '1' & x"02";
tmp(218) := 								RET & "00" & '0' & x"00";
tmp(219) := 										LDI & "00" & '0' & x"01";
tmp(220) := 										STA & "00" & '0' & x"16";
tmp(221) := 										STA & "00" & '1' & x"02";
tmp(222) := 										RET & "00" & '0' & x"00";
tmp(223) := 	STA & "10" & '1' & x"20";
tmp(224) := 	STA & "11" & '1' & x"21";
tmp(225) := 	LDA & "01" & '0' & x"00";
tmp(226) := 	STA & "01" & '1' & x"22";
tmp(227) := 	LDA & "01" & '0' & x"01";
tmp(228) := 	STA & "01" & '1' & x"23";
tmp(229) := 	LDA & "01" & '0' & x"02";
tmp(230) := 	STA & "01" & '1' & x"24";
tmp(231) := 	LDA & "01" & '0' & x"03";
tmp(232) := 	STA & "01" & '1' & x"25";
tmp(233) := 	RET & "00" & '0' & x"00";
tmp(234) := 	CEQ & "10" & '0' & x"1E";
tmp(235) := 	JEQ & "00" & '0' & x"ED";
tmp(236) := 	RET & "00" & '0' & x"00";
tmp(237) := 		CEQ & "11" & '0' & x"1F";
tmp(238) := 		JEQ & "00" & '0' & x"F0";
tmp(239) := 		RET & "00" & '0' & x"00";
tmp(240) := 			LDA & "00" & '0' & x"00";
tmp(241) := 			CEQ & "00" & '0' & x"20";
tmp(242) := 			JEQ & "00" & '0' & x"F4";
tmp(243) := 			RET & "00" & '0' & x"00";
tmp(244) := 				LDA & "00" & '0' & x"01";
tmp(245) := 				CEQ & "00" & '0' & x"21";
tmp(246) := 				JEQ & "00" & '0' & x"F8";
tmp(247) := 				RET & "00" & '0' & x"00";
tmp(248) := 					LDA & "00" & '0' & x"02";
tmp(249) := 					CEQ & "00" & '0' & x"22";
tmp(250) := 					JEQ & "00" & '0' & x"FC";
tmp(251) := 					RET & "00" & '0' & x"00";
tmp(252) := 						LDA & "00" & '0' & x"03";
tmp(253) := 						CEQ & "00" & '0' & x"23";
tmp(254) := 						JEQ & "00" & '1' & x"00";
tmp(255) := 						RET & "00" & '0' & x"00";
tmp(256) := 							LDI & "00" & '0' & x"00";
tmp(257) := 							STA & "00" & '0' & x"14";
tmp(258) := 							LDI & "00" & '0' & x"01";
tmp(259) := 							STA & "00" & '1' & x"01";
tmp(260) := 							LDI & "00" & '0' & x"00";
tmp(261) := 							RET & "00" & '0' & x"00";

        
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;