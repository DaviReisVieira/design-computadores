LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY logicaDesvio IS

  PORT (
    JLT, JMP, JEQ, JSR, RET : IN STD_LOGIC;
    FLAG_EQ : IN STD_LOGIC;
    FLAG_LESS : IN STD_LOGIC;
    Sel : OUT std_logic_vector(1 downto 0)
  );
END ENTITY;
ARCHITECTURE arch_name OF logicaDesvio IS

-- CONTROLA A PORTA DO MUX 4X1, CUJA SAÍDA É O ENDEREÇO DA PRÓXIMA INSTRUÇÃO
-- 00: Próximo PC
-- 01: Endereço Imediato
-- 02: Endereço Retorno
-- 03: Aberto.

BEGIN

Sel(1) <= NOT JMP AND RET AND NOT JSR AND NOT JEQ AND NOT JLT;

Sel(0) <= (JMP AND NOT RET AND NOT JSR AND NOT JEQ AND NOT JLT) OR 
				  (NOT JMP AND NOT RET AND NOT JSR AND JEQ AND NOT JLT AND FLAG_EQ AND NOT FLAG_LESS) OR 
				  (NOT JMP AND NOT RET AND NOT JSR AND NOT JEQ AND JLT AND NOT FLAG_EQ AND FLAG_LESS) OR 
				  (NOT JMP AND NOT RET AND JSR AND NOT JEQ AND NOT JLT);

END ARCHITECTURE;