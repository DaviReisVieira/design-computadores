library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 15;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
  constant RET  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin      

  tmp(0) :=     LDI & "00" & '0' & x"00";
tmp(1) := 	LDI & "01" & '0' & x"00";
tmp(2) := 	LDI & "10" & '0' & x"00";
tmp(3) := 	LDI & "11" & '0' & x"00";
tmp(4) := 	STA & "00" & '1' & x"20";
tmp(5) := 	STA & "00" & '1' & x"21";
tmp(6) := 	STA & "00" & '1' & x"22";
tmp(7) := 	STA & "00" & '1' & x"23";
tmp(8) := 	STA & "00" & '1' & x"24";
tmp(9) := 	STA & "00" & '1' & x"25";
tmp(10) := 	STA & "00" & '1' & x"00";
tmp(11) := 	STA & "00" & '1' & x"01";
tmp(12) := 	STA & "00" & '1' & x"02";
tmp(13) := 	STA & "00" & '0' & x"00";
tmp(14) := 	STA & "00" & '0' & x"01";
tmp(15) := 	STA & "00" & '0' & x"02";
tmp(16) := 	STA & "00" & '0' & x"03";
tmp(17) := 	LDI & "00" & '0' & x"09";
tmp(18) := 	STA & "00" & '0' & x"1E";
tmp(19) := 	STA & "00" & '0' & x"1F";
tmp(20) := 	STA & "00" & '0' & x"20";
tmp(21) := 	STA & "00" & '0' & x"21";
tmp(22) := 	STA & "00" & '0' & x"22";
tmp(23) := 	STA & "00" & '0' & x"23";
tmp(24) := 	LDI & "00" & '0' & x"00";
tmp(25) := 	STA & "00" & '0' & x"0A";
tmp(26) := 	LDI & "00" & '0' & x"01";
tmp(27) := 	STA & "00" & '0' & x"0B";
tmp(28) := 	LDI & "00" & '0' & x"0A";
tmp(29) := 	STA & "00" & '0' & x"0C";
tmp(30) := 	LDI & "00" & '0' & x"01";
tmp(31) := 	STA & "00" & '0' & x"14";
tmp(32) := 	LDI & "00" & '0' & x"00";
tmp(33) := 	STA & "00" & '1' & x"FE";
tmp(34) := 	STA & "00" & '1' & x"FC";
tmp(35) := 	STA & "00" & '1' & x"FD";
tmp(36) := 	LDA & "01" & '1' & x"65";
tmp(37) := 	CEQ & "01" & '0' & x"0A";
tmp(38) := 	JSR & "00" & '0' & x"B7";
tmp(39) := 	JEQ & "00" & '0' & x"2E";
tmp(40) := 	JSR & "00" & '0' & x"C2";
tmp(41) := 	JSR & "00" & '0' & x"86";
tmp(42) := 	LDA & "01" & '1' & x"64";
tmp(43) := 	CEQ & "01" & '0' & x"0A";
tmp(44) := 	JEQ & "00" & '0' & x"2E";
tmp(45) := 	JSR & "00" & '0' & x"74";
tmp(46) := 			LDA & "01" & '1' & x"61";
tmp(47) := 			CEQ & "01" & '0' & x"0A";
tmp(48) := 			JEQ & "00" & '0' & x"72";
tmp(49) := 			STA & "00" & '1' & x"FE";
tmp(50) := 				LDI & "00" & '0' & x"01";
tmp(51) := 				STA & "00" & '1' & x"00";
tmp(52) := 					LDA & "00" & '1' & x"40";
tmp(53) := 					STA & "00" & '1' & x"20";
tmp(54) := 					LDA & "01" & '1' & x"61";
tmp(55) := 					CEQ & "01" & '0' & x"0A";
tmp(56) := 					JEQ & "00" & '0' & x"34";
tmp(57) := 					STA & "00" & '1' & x"FE";
tmp(58) := 					STA & "00" & '0' & x"1E";
tmp(59) := 				LDI & "00" & '0' & x"02";
tmp(60) := 				STA & "00" & '1' & x"00";
tmp(61) := 					LDA & "00" & '1' & x"40";
tmp(62) := 					STA & "00" & '1' & x"21";
tmp(63) := 					LDA & "01" & '1' & x"61";
tmp(64) := 					CEQ & "01" & '0' & x"0A";
tmp(65) := 					JEQ & "00" & '0' & x"3D";
tmp(66) := 					STA & "00" & '1' & x"FE";
tmp(67) := 					STA & "00" & '0' & x"1F";
tmp(68) := 				LDI & "00" & '0' & x"04";
tmp(69) := 				STA & "00" & '1' & x"00";
tmp(70) := 					LDA & "00" & '1' & x"40";
tmp(71) := 					STA & "00" & '1' & x"22";
tmp(72) := 					LDA & "01" & '1' & x"61";
tmp(73) := 					CEQ & "01" & '0' & x"0A";
tmp(74) := 					JEQ & "00" & '0' & x"46";
tmp(75) := 					STA & "00" & '1' & x"FE";
tmp(76) := 					STA & "00" & '0' & x"20";
tmp(77) := 				LDI & "00" & '0' & x"08";
tmp(78) := 				STA & "00" & '1' & x"00";
tmp(79) := 					LDA & "00" & '1' & x"40";
tmp(80) := 					STA & "00" & '1' & x"23";
tmp(81) := 					LDA & "01" & '1' & x"61";
tmp(82) := 					CEQ & "01" & '0' & x"0A";
tmp(83) := 					JEQ & "00" & '0' & x"4F";
tmp(84) := 					STA & "00" & '1' & x"FE";
tmp(85) := 					STA & "00" & '0' & x"21";
tmp(86) := 				LDI & "00" & '0' & x"10";
tmp(87) := 				STA & "00" & '1' & x"00";
tmp(88) := 					LDA & "00" & '1' & x"40";
tmp(89) := 					STA & "00" & '1' & x"24";
tmp(90) := 					LDA & "01" & '1' & x"61";
tmp(91) := 					CEQ & "01" & '0' & x"0A";
tmp(92) := 					JEQ & "00" & '0' & x"58";
tmp(93) := 					STA & "00" & '1' & x"FE";
tmp(94) := 					STA & "00" & '0' & x"22";
tmp(95) := 				LDI & "00" & '0' & x"20";
tmp(96) := 				STA & "00" & '1' & x"00";
tmp(97) := 					LDA & "00" & '1' & x"40";
tmp(98) := 					STA & "00" & '1' & x"25";
tmp(99) := 					LDA & "01" & '1' & x"61";
tmp(100) := 					CEQ & "01" & '0' & x"0A";
tmp(101) := 					JEQ & "00" & '0' & x"61";
tmp(102) := 					STA & "00" & '1' & x"FE";
tmp(103) := 					STA & "00" & '0' & x"23";
tmp(104) := 					LDI & "00" & '0' & x"00";
tmp(105) := 					LDI & "01" & '0' & x"00";
tmp(106) := 					STA & "00" & '1' & x"00";
tmp(107) := 					LDI & "00" & '0' & x"00";
tmp(108) := 					STA & "00" & '1' & x"20";
tmp(109) := 					STA & "00" & '1' & x"21";
tmp(110) := 					STA & "00" & '1' & x"22";
tmp(111) := 					STA & "00" & '1' & x"23";
tmp(112) := 					STA & "00" & '1' & x"24";
tmp(113) := 					STA & "00" & '1' & x"25";
tmp(114) := 				NOP & "00" & '0' & x"00";
tmp(115) := JMP  & "00" & '0' & x"24";
tmp(116) := 	STA & "00" & '1' & x"FD";
tmp(117) := 	LDI & "10" & '0' & x"00";
tmp(118) := 	STA & "10" & '0' & x"00";
tmp(119) := 	STA & "10" & '0' & x"01";
tmp(120) := 	STA & "10" & '0' & x"02";
tmp(121) := 	STA & "10" & '0' & x"03";
tmp(122) := 	STA & "10" & '1' & x"20";
tmp(123) := 	STA & "10" & '1' & x"21";
tmp(124) := 	STA & "10" & '1' & x"22";
tmp(125) := 	STA & "10" & '1' & x"23";
tmp(126) := 	STA & "10" & '1' & x"24";
tmp(127) := 	STA & "10" & '1' & x"25";
tmp(128) := 	STA & "10" & '1' & x"01";
tmp(129) := 	STA & "10" & '1' & x"02";
tmp(130) := 	LDI & "11" & '0' & x"01";
tmp(131) := 	STA & "11" & '0' & x"14";
tmp(132) := 	LDI & "11" & '0' & x"00";
tmp(133) := 	RET & "00" & '0' & x"00";
tmp(134) := 	STA & "00" & '1' & x"FC";
tmp(135) := 	LDA & "01" & '0' & x"14";
tmp(136) := 	CEQ & "01" & '0' & x"0B";
tmp(137) := 	JEQ & "00" & '0' & x"8B";
tmp(138) := 	RET & "00" & '0' & x"00";
tmp(139) := 		SOMA & "10" & '0' & x"0B";
tmp(140) := 		CEQ & "10" & '0' & x"0C";
tmp(141) := 		JEQ & "00" & '0' & x"8F";
tmp(142) := 		RET & "00" & '0' & x"00";
tmp(143) := 			SOMA & "11" & '0' & x"0B";
tmp(144) := 			CEQ & "11" & '0' & x"0C";
tmp(145) := 			LDI & "10" & '0' & x"00";
tmp(146) := 			JEQ & "00" & '0' & x"94";
tmp(147) := 			RET & "00" & '0' & x"00";
tmp(148) := 				LDI & "00" & '0' & x"01";
tmp(149) := 				SOMA & "00" & '0' & x"00";
tmp(150) := 				LDI & "11" & '0' & x"00";
tmp(151) := 				CEQ & "00" & '0' & x"0C";
tmp(152) := 				JEQ & "00" & '0' & x"9B";
tmp(153) := 				STA & "00" & '0' & x"00";
tmp(154) := 				RET & "00" & '0' & x"00";
tmp(155) := 					LDI & "00" & '0' & x"00";
tmp(156) := 					STA & "00" & '0' & x"00";
tmp(157) := 					LDI & "00" & '0' & x"01";
tmp(158) := 					SOMA & "00" & '0' & x"01";
tmp(159) := 					CEQ & "00" & '0' & x"0C";
tmp(160) := 					JEQ & "00" & '0' & x"A3";
tmp(161) := 					STA & "00" & '0' & x"01";
tmp(162) := 					RET & "00" & '0' & x"00";
tmp(163) := 						LDI & "00" & '0' & x"00";
tmp(164) := 						STA & "00" & '0' & x"01";
tmp(165) := 						LDI & "00" & '0' & x"01";
tmp(166) := 						SOMA & "00" & '0' & x"02";
tmp(167) := 						CEQ & "00" & '0' & x"0C";
tmp(168) := 						JEQ & "00" & '0' & x"AB";
tmp(169) := 						STA & "00" & '0' & x"02";
tmp(170) := 						RET & "00" & '0' & x"00";
tmp(171) := 							LDI & "00" & '0' & x"00";
tmp(172) := 							STA & "00" & '0' & x"02";
tmp(173) := 							LDI & "00" & '0' & x"01";
tmp(174) := 							SOMA & "00" & '0' & x"03";
tmp(175) := 							CEQ & "00" & '0' & x"0C";
tmp(176) := 							JEQ & "00" & '0' & x"B2";
tmp(177) := 							RET & "00" & '0' & x"00";
tmp(178) := 								LDI & "00" & '0' & x"01";
tmp(179) := 								STA & "00" & '1' & x"02";
tmp(180) := 								LDI & "00" & '0' & x"00";
tmp(181) := 								STA & "00" & '0' & x"14";
tmp(182) := 								RET & "00" & '0' & x"00";
tmp(183) := 	STA & "10" & '1' & x"20";
tmp(184) := 	STA & "11" & '1' & x"21";
tmp(185) := 	LDA & "01" & '0' & x"00";
tmp(186) := 	STA & "01" & '1' & x"22";
tmp(187) := 	LDA & "01" & '0' & x"01";
tmp(188) := 	STA & "01" & '1' & x"23";
tmp(189) := 	LDA & "01" & '0' & x"02";
tmp(190) := 	STA & "01" & '1' & x"24";
tmp(191) := 	LDA & "01" & '0' & x"03";
tmp(192) := 	STA & "01" & '1' & x"25";
tmp(193) := 	RET & "00" & '0' & x"00";
tmp(194) := 	CEQ & "10" & '0' & x"1E";
tmp(195) := 	JEQ & "00" & '0' & x"C5";
tmp(196) := 	RET & "00" & '0' & x"00";
tmp(197) := 		CEQ & "11" & '0' & x"1F";
tmp(198) := 		JEQ & "00" & '0' & x"C8";
tmp(199) := 		RET & "00" & '0' & x"00";
tmp(200) := 			LDA & "00" & '0' & x"00";
tmp(201) := 			CEQ & "00" & '0' & x"20";
tmp(202) := 			JEQ & "00" & '0' & x"CC";
tmp(203) := 			RET & "00" & '0' & x"00";
tmp(204) := 				LDA & "00" & '0' & x"01";
tmp(205) := 				CEQ & "00" & '0' & x"21";
tmp(206) := 				JEQ & "00" & '0' & x"D0";
tmp(207) := 				RET & "00" & '0' & x"00";
tmp(208) := 					LDA & "00" & '0' & x"02";
tmp(209) := 					CEQ & "00" & '0' & x"22";
tmp(210) := 					JEQ & "00" & '0' & x"D4";
tmp(211) := 					RET & "00" & '0' & x"00";
tmp(212) := 						LDA & "00" & '0' & x"03";
tmp(213) := 						CEQ & "00" & '0' & x"23";
tmp(214) := 						JEQ & "00" & '0' & x"D8";
tmp(215) := 						RET & "00" & '0' & x"00";
tmp(216) := 							LDI & "00" & '0' & x"00";
tmp(217) := 							STA & "00" & '0' & x"14";
tmp(218) := 							LDI & "00" & '0' & x"01";
tmp(219) := 							STA & "00" & '1' & x"01";
tmp(220) := 							LDI & "00" & '0' & x"00";
tmp(221) := 							RET & "00" & '0' & x"00";

        
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;