library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 15;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
  constant RET  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
  constant CLT  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1011";
  constant JLT  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1100";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin      

  tmp(0) :=     LDI & "00" & '0' & x"00";
  tmp(1) := 	LDI & "01" & '0' & x"00";
  tmp(2) := 	LDI & "10" & '0' & x"00";
  tmp(3) := 	LDI & "11" & '0' & x"00";
  tmp(4) := 	STA & "00" & '1' & x"00";
  tmp(5) := 	STA & "00" & '1' & x"01";
  tmp(6) := 	STA & "00" & '1' & x"02";
  tmp(7) := 	STA & "00" & '0' & x"00";
  tmp(8) := 	STA & "00" & '0' & x"01";
  tmp(9) := 	STA & "00" & '0' & x"02";
  tmp(10) := 	STA & "00" & '0' & x"03";
  tmp(11) := 	LDI & "00" & '0' & x"09";
  tmp(12) := 	STA & "00" & '0' & x"1E";
  tmp(13) := 	STA & "00" & '0' & x"1F";
  tmp(14) := 	STA & "00" & '0' & x"20";
  tmp(15) := 	STA & "00" & '0' & x"21";
  tmp(16) := 	STA & "00" & '0' & x"22";
  tmp(17) := 	STA & "00" & '0' & x"23";
  tmp(18) := 	LDI & "00" & '0' & x"00";
  tmp(19) := 	STA & "00" & '0' & x"0A";
  tmp(20) := 	LDI & "00" & '0' & x"01";
  tmp(21) := 	STA & "00" & '0' & x"0B";
  tmp(22) := 	LDI & "00" & '0' & x"0A";
  tmp(23) := 	STA & "00" & '0' & x"0C";
  tmp(24) := 	LDI & "00" & '0' & x"06";
  tmp(25) := 	STA & "00" & '0' & x"0D";
  tmp(26) := 	LDI & "00" & '0' & x"04";
  tmp(27) := 	STA & "00" & '0' & x"0E";
  tmp(28) := 	LDI & "00" & '0' & x"02";
  tmp(29) := 	STA & "00" & '0' & x"0F";
  tmp(30) := 	LDI & "00" & '0' & x"01";
  tmp(31) := 	STA & "00" & '0' & x"14";
  tmp(32) := 	LDI & "00" & '0' & x"01";
  tmp(33) := 	STA & "00" & '0' & x"15";
  tmp(34) := 	LDI & "00" & '0' & x"00";
  tmp(35) := 	STA & "00" & '0' & x"16";
  tmp(36) := 	LDI & "00" & '0' & x"01";
  tmp(37) := 	STA & "00" & '0' & x"17";
  tmp(38) := 	LDI & "00" & '0' & x"00";
  tmp(39) := 	STA & "00" & '1' & x"FE";
  tmp(40) := 	STA & "00" & '1' & x"FC";
  tmp(41) := 	STA & "00" & '1' & x"FD";
  tmp(42) := 	LDA & "01" & '1' & x"65";
  tmp(43) := 	CEQ & "01" & '0' & x"0A";
  tmp(44) := 	JSR & "00" & '1' & x"CF";
  tmp(45) := 	JEQ & "00" & '0' & x"34";
  tmp(46) := 	JSR & "00" & '1' & x"DE";
  tmp(47) := 	JSR & "00" & '1' & x"82";
  tmp(48) := 	LDA & "01" & '1' & x"64";
  tmp(49) := 	CEQ & "01" & '0' & x"0A";
  tmp(50) := 	JEQ & "00" & '0' & x"34";
  tmp(51) := 	JSR & "00" & '1' & x"78";
  tmp(52) := 			LDA & "01" & '1' & x"61";
  tmp(53) := 			CEQ & "01" & '0' & x"0A";
  tmp(54) := 			JEQ & "00" & '0' & x"3B";
  tmp(55) := 			STA & "00" & '1' & x"FE";
  tmp(56) := 			LDI & "00" & '0' & x"00";
  tmp(57) := 			STA & "00" & '0' & x"17";
  tmp(58) := 			JSR & "00" & '0' & x"A0";
  tmp(59) := 				STA & "00" & '1' & x"FE";
  tmp(60) := 				LDA & "01" & '1' & x"60";
  tmp(61) := 				CEQ & "01" & '0' & x"0A";
  tmp(62) := 				JEQ & "00" & '0' & x"42";
  tmp(63) := 				LDI & "00" & '0' & x"01";
  tmp(64) := 				STA & "00" & '0' & x"17";
  tmp(65) := 				JSR & "00" & '0' & x"A0";
  tmp(66) := 					LDA & "01" & '1' & x"62";
  tmp(67) := 					CEQ & "01" & '0' & x"0A";
  tmp(68) := 					JEQ & "00" & '0' & x"46";
  tmp(69) := 					JSR & "00" & '0' & x"48";
  tmp(70) := 						NOP & "00" & '0' & x"00";
  tmp(71) := JMP  & "00" & '0' & x"2A";
  tmp(72) := 	STA & "00" & '1' & x"FB";
  tmp(73) := 	LDA & "00" & '0' & x"15";
  tmp(74) := 	CEQ & "00" & '0' & x"0A";
  tmp(75) := 	JEQ & "00" & '0' & x"86";
  tmp(76) := 	LDI & "00" & '0' & x"00";
  tmp(77) := 	STA & "00" & '0' & x"15";
  tmp(78) := 		LDA & "00" & '0' & x"03";
  tmp(79) := 		CEQ & "00" & '0' & x"0B";
  tmp(80) := 		JEQ & "00" & '0' & x"54";
  tmp(81) := 		CEQ & "00" & '0' & x"0F";
  tmp(82) := 		JEQ & "00" & '0' & x"62";
  tmp(83) := 		RET & "00" & '0' & x"00";
  tmp(84) := 			LDI & "00" & '0' & x"01";
  tmp(85) := 			CLT & "00" & '0' & x"02";
  tmp(86) := 			JLT & "00" & '0' & x"58";
  tmp(87) := 			RET & "00" & '0' & x"00";
  tmp(88) := 				LDA & "00" & '0' & x"02";
  tmp(89) := 				SUB & "00" & '0' & x"0F";
  tmp(90) := 				STA & "00" & '0' & x"02";
  tmp(91) := 				STA & "00" & '0' & x"22";
  tmp(92) := 				LDI & "00" & '0' & x"00";
  tmp(93) := 				STA & "00" & '0' & x"03";
  tmp(94) := 				STA & "00" & '0' & x"23";
  tmp(95) := 				LDI & "00" & '0' & x"01";
  tmp(96) := 				STA & "00" & '0' & x"16";
  tmp(97) := 				RET & "00" & '0' & x"00";
  tmp(98) := 			LDI & "00" & '0' & x"01";
  tmp(99) := 			STA & "00" & '0' & x"16";
  tmp(100) := 			LDA & "00" & '0' & x"02";
  tmp(101) := 			CEQ & "00" & '0' & x"0A";
  tmp(102) := 			JEQ & "00" & '0' & x"6C";
  tmp(103) := 			CEQ & "00" & '0' & x"0B";
  tmp(104) := 			JEQ & "00" & '0' & x"72";
  tmp(105) := 			CEQ & "00" & '0' & x"0F";
  tmp(106) := 			JEQ & "00" & '0' & x"79";
  tmp(107) := 			JMP & "00" & '0' & x"80";
  tmp(108) := 				LDI & "01" & '0' & x"08";
  tmp(109) := 				STA & "01" & '0' & x"02";
  tmp(110) := 				STA & "01" & '0' & x"22";
  tmp(111) := 				STA & "00" & '0' & x"03";
  tmp(112) := 				STA & "00" & '0' & x"23";
  tmp(113) := 				RET & "00" & '0' & x"00";
  tmp(114) := 				LDI & "01" & '0' & x"09";
  tmp(115) := 				STA & "01" & '0' & x"02";
  tmp(116) := 				STA & "01" & '0' & x"22";
  tmp(117) := 				LDI & "00" & '0' & x"00";
  tmp(118) := 				STA & "00" & '0' & x"03";
  tmp(119) := 				STA & "00" & '0' & x"23";
  tmp(120) := 				RET & "00" & '0' & x"00";
  tmp(121) := 				LDI & "00" & '0' & x"00";
  tmp(122) := 				STA & "00" & '0' & x"02";
  tmp(123) := 				STA & "00" & '0' & x"22";
  tmp(124) := 				LDI & "01" & '0' & x"01";
  tmp(125) := 				STA & "01" & '0' & x"03";
  tmp(126) := 				STA & "01" & '0' & x"23";
  tmp(127) := 				RET & "00" & '0' & x"00";
  tmp(128) := 				LDI & "01" & '0' & x"01";
  tmp(129) := 				STA & "01" & '0' & x"02";
  tmp(130) := 				STA & "01" & '0' & x"22";
  tmp(131) := 				STA & "01" & '0' & x"03";
  tmp(132) := 				STA & "01" & '0' & x"23";
  tmp(133) := 				RET & "00" & '0' & x"00";
  tmp(134) := 		LDI & "00" & '0' & x"01";
  tmp(135) := 		STA & "00" & '0' & x"15";
  tmp(136) := 		LDA & "00" & '0' & x"16";
  tmp(137) := 		CEQ & "00" & '0' & x"0A";
  tmp(138) := 		JEQ & "00" & '0' & x"9D";
  tmp(139) := 		LDA & "00" & '0' & x"02";
  tmp(140) := 		SOMA & "00" & '0' & x"0F";
  tmp(141) := 		STA & "00" & '0' & x"02";
  tmp(142) := 		LDI & "00" & '0' & x"09";
  tmp(143) := 		CLT & "00" & '0' & x"02";
  tmp(144) := 		JLT & "00" & '0' & x"92";
  tmp(145) := 		JMP & "00" & '0' & x"99";
  tmp(146) := 			LDA & "00" & '0' & x"02";
  tmp(147) := 			SUB & "00" & '0' & x"0C";
  tmp(148) := 			STA & "00" & '0' & x"02";
  tmp(149) := 			STA & "00" & '0' & x"22";
  tmp(150) := 			LDA & "00" & '0' & x"03";
  tmp(151) := 			SOMA & "00" & '0' & x"0B";
  tmp(152) := 			STA & "00" & '0' & x"03";
  tmp(153) := 			LDA & "00" & '0' & x"03";
  tmp(154) := 			SOMA & "00" & '0' & x"0B";
  tmp(155) := 			STA & "00" & '0' & x"03";
  tmp(156) := 			STA & "00" & '0' & x"23";
  tmp(157) := 			LDI & "00" & '0' & x"00";
  tmp(158) := 			STA & "00" & '0' & x"16";
  tmp(159) := 			RET & "00" & '0' & x"00";
  tmp(160) := 	LDI & "00" & '0' & x"00";
  tmp(161) := 	STA & "00" & '1' & x"20";
  tmp(162) := 	STA & "00" & '1' & x"21";
  tmp(163) := 	STA & "00" & '1' & x"22";
  tmp(164) := 	STA & "00" & '1' & x"23";
  tmp(165) := 	STA & "00" & '1' & x"24";
  tmp(166) := 	STA & "00" & '1' & x"25";
  tmp(167) := 		STA & "00" & '1' & x"FE";
  tmp(168) := 		STA & "00" & '1' & x"FF";
  tmp(169) := 		LDI & "00" & '0' & x"01";
  tmp(170) := 		STA & "00" & '1' & x"02";
  tmp(171) := 			LDA & "00" & '1' & x"40";
  tmp(172) := 			LDA & "01" & '0' & x"15";
  tmp(173) := 			CEQ & "01" & '0' & x"0A";
  tmp(174) := 			JEQ & "00" & '0' & x"C0";
  tmp(175) := 			LDI & "01" & '0' & x"02";
  tmp(176) := 			CLT & "01" & '1' & x"40";
  tmp(177) := 			JLT & "00" & '0' & x"B3";
  tmp(178) := 			JMP & "00" & '0' & x"B4";
  tmp(179) := 				LDI & "00" & '0' & x"02";
  tmp(180) := 				STA & "00" & '1' & x"25";
  tmp(181) := 				LDA & "01" & '1' & x"60";
  tmp(182) := 				CEQ & "01" & '0' & x"0A";
  tmp(183) := 				JEQ & "00" & '0' & x"AB";
  tmp(184) := 				STA & "00" & '1' & x"FF";
  tmp(185) := 				LDA & "01" & '0' & x"17";
  tmp(186) := 				CEQ & "01" & '0' & x"0B";
  tmp(187) := 				JEQ & "00" & '0' & x"BE";
  tmp(188) := 				STA & "00" & '0' & x"23";
  tmp(189) := 				JMP & "00" & '0' & x"D0";
  tmp(190) := 					STA & "00" & '0' & x"03";
  tmp(191) := 					JMP & "00" & '0' & x"D0";
  tmp(192) := 				LDI & "01" & '0' & x"01";
  tmp(193) := 				CLT & "01" & '1' & x"40";
  tmp(194) := 				JLT & "00" & '0' & x"C4";
  tmp(195) := 				JMP & "00" & '0' & x"C5";
  tmp(196) := 					LDI & "00" & '0' & x"01";
  tmp(197) := 					STA & "00" & '1' & x"25";
  tmp(198) := 					LDA & "01" & '1' & x"60";
  tmp(199) := 					CEQ & "01" & '0' & x"0A";
  tmp(200) := 					JEQ & "00" & '0' & x"AB";
  tmp(201) := 					STA & "00" & '1' & x"FF";
  tmp(202) := 					LDA & "01" & '0' & x"17";
  tmp(203) := 					CEQ & "01" & '0' & x"0B";
  tmp(204) := 					JEQ & "00" & '0' & x"CF";
  tmp(205) := 					STA & "00" & '0' & x"23";
  tmp(206) := 					JMP & "00" & '0' & x"D0";
  tmp(207) := 						STA & "00" & '0' & x"03";
  tmp(208) := 		STA & "00" & '1' & x"FF";
  tmp(209) := 		LDI & "00" & '0' & x"01";
  tmp(210) := 		STA & "00" & '1' & x"01";
  tmp(211) := 			LDA & "00" & '1' & x"40";
  tmp(212) := 			LDA & "01" & '0' & x"15";
  tmp(213) := 			CEQ & "01" & '0' & x"0A";
  tmp(214) := 			JEQ & "00" & '0' & x"FC";
  tmp(215) := 			LDI & "01" & '0' & x"02";
  tmp(216) := 			CEQ & "01" & '0' & x"03";
  tmp(217) := 			JEQ & "00" & '0' & x"EB";
  tmp(218) := 			LDI & "01" & '0' & x"0A";
  tmp(219) := 			CLT & "01" & '1' & x"40";
  tmp(220) := 			JLT & "00" & '0' & x"DE";
  tmp(221) := 			JMP & "00" & '0' & x"DF";
  tmp(222) := 				LDI & "00" & '0' & x"09";
  tmp(223) := 				STA & "00" & '1' & x"24";
  tmp(224) := 				LDA & "01" & '1' & x"60";
  tmp(225) := 				CEQ & "01" & '0' & x"0A";
  tmp(226) := 				JEQ & "00" & '0' & x"D3";
  tmp(227) := 				STA & "00" & '1' & x"FF";
  tmp(228) := 				LDA & "01" & '0' & x"17";
  tmp(229) := 				CEQ & "01" & '0' & x"0B";
  tmp(230) := 				JEQ & "00" & '0' & x"E9";
  tmp(231) := 				STA & "00" & '0' & x"22";
  tmp(232) := 				JMP & "00" & '1' & x"20";
  tmp(233) := 					STA & "00" & '0' & x"02";
  tmp(234) := 					JMP & "00" & '1' & x"20";
  tmp(235) := 				LDI & "01" & '0' & x"03";
  tmp(236) := 				CLT & "01" & '1' & x"40";
  tmp(237) := 				JLT & "00" & '0' & x"EF";
  tmp(238) := 				JMP & "00" & '0' & x"F0";
  tmp(239) := 					LDI & "00" & '0' & x"03";
  tmp(240) := 					STA & "00" & '1' & x"24";
  tmp(241) := 					LDA & "01" & '1' & x"60";
  tmp(242) := 					CEQ & "01" & '0' & x"0A";
  tmp(243) := 					JEQ & "00" & '0' & x"D3";
  tmp(244) := 					STA & "00" & '1' & x"FF";
  tmp(245) := 					LDA & "01" & '0' & x"17";
  tmp(246) := 					CEQ & "01" & '0' & x"0B";
  tmp(247) := 					JEQ & "00" & '0' & x"FA";
  tmp(248) := 					STA & "00" & '0' & x"22";
  tmp(249) := 					JMP & "00" & '1' & x"20";
  tmp(250) := 						STA & "00" & '0' & x"02";
  tmp(251) := 						JMP & "00" & '1' & x"20";
  tmp(252) := 				LDI & "01" & '0' & x"01";
  tmp(253) := 				CEQ & "01" & '0' & x"03";
  tmp(254) := 				JEQ & "00" & '1' & x"10";
  tmp(255) := 				LDI & "01" & '0' & x"0A";
  tmp(256) := 				CLT & "01" & '1' & x"40";
  tmp(257) := 				JLT & "00" & '1' & x"03";
  tmp(258) := 				JMP & "00" & '1' & x"04";
  tmp(259) := 					LDI & "00" & '0' & x"09";
  tmp(260) := 					STA & "00" & '1' & x"24";
  tmp(261) := 					LDA & "01" & '1' & x"60";
  tmp(262) := 					CEQ & "01" & '0' & x"0A";
  tmp(263) := 					JEQ & "00" & '0' & x"D3";
  tmp(264) := 					STA & "00" & '1' & x"FF";
  tmp(265) := 					LDA & "01" & '0' & x"17";
  tmp(266) := 					CEQ & "01" & '0' & x"0B";
  tmp(267) := 					JEQ & "00" & '1' & x"0E";
  tmp(268) := 					STA & "00" & '0' & x"22";
  tmp(269) := 					JMP & "00" & '1' & x"20";
  tmp(270) := 						STA & "00" & '0' & x"02";
  tmp(271) := 						JMP & "00" & '1' & x"20";
  tmp(272) := 					LDI & "01" & '0' & x"02";
  tmp(273) := 					CLT & "01" & '1' & x"40";
  tmp(274) := 					JLT & "00" & '1' & x"14";
  tmp(275) := 					JMP & "00" & '1' & x"15";
  tmp(276) := 						LDI & "00" & '0' & x"01";
  tmp(277) := 						STA & "00" & '1' & x"24";
  tmp(278) := 						LDA & "01" & '1' & x"60";
  tmp(279) := 						CEQ & "01" & '0' & x"0A";
  tmp(280) := 						JEQ & "00" & '0' & x"D3";
  tmp(281) := 						STA & "00" & '1' & x"FF";
  tmp(282) := 						LDA & "01" & '0' & x"17";
  tmp(283) := 						CEQ & "01" & '0' & x"0B";
  tmp(284) := 						JEQ & "00" & '1' & x"1F";
  tmp(285) := 						STA & "00" & '0' & x"22";
  tmp(286) := 						JMP & "00" & '1' & x"20";
  tmp(287) := 							STA & "00" & '0' & x"02";
  tmp(288) := 		STA & "00" & '1' & x"FF";
  tmp(289) := 		LDI & "00" & '0' & x"80";
  tmp(290) := 		STA & "00" & '1' & x"00";
  tmp(291) := 			LDA & "00" & '1' & x"40";
  tmp(292) := 			LDI & "01" & '0' & x"06";
  tmp(293) := 			CLT & "01" & '1' & x"40";
  tmp(294) := 			JLT & "00" & '1' & x"28";
  tmp(295) := 			JMP & "00" & '1' & x"29";
  tmp(296) := 				LDI & "00" & '0' & x"05";
  tmp(297) := 				STA & "00" & '1' & x"23";
  tmp(298) := 				LDA & "01" & '1' & x"60";
  tmp(299) := 				CEQ & "01" & '0' & x"0A";
  tmp(300) := 				JEQ & "00" & '1' & x"23";
  tmp(301) := 				STA & "00" & '1' & x"FF";
  tmp(302) := 				LDA & "01" & '0' & x"17";
  tmp(303) := 				CEQ & "01" & '0' & x"0B";
  tmp(304) := 				JEQ & "00" & '1' & x"33";
  tmp(305) := 				STA & "00" & '0' & x"21";
  tmp(306) := 				JMP & "00" & '1' & x"34";
  tmp(307) := 					STA & "00" & '0' & x"01";
  tmp(308) := 		STA & "00" & '1' & x"FF";
  tmp(309) := 		LDI & "00" & '0' & x"C0";
  tmp(310) := 		STA & "00" & '1' & x"00";
  tmp(311) := 			LDA & "00" & '1' & x"40";
  tmp(312) := 			LDI & "01" & '0' & x"0A";
  tmp(313) := 			CLT & "01" & '1' & x"40";
  tmp(314) := 			JLT & "00" & '1' & x"3C";
  tmp(315) := 			JMP & "00" & '1' & x"3D";
  tmp(316) := 				LDI & "00" & '0' & x"09";
  tmp(317) := 				STA & "00" & '1' & x"22";
  tmp(318) := 				LDA & "01" & '1' & x"60";
  tmp(319) := 				CEQ & "01" & '0' & x"0A";
  tmp(320) := 				JEQ & "00" & '1' & x"37";
  tmp(321) := 				STA & "00" & '1' & x"FF";
  tmp(322) := 				LDA & "01" & '0' & x"17";
  tmp(323) := 				CEQ & "01" & '0' & x"0B";
  tmp(324) := 				JEQ & "00" & '1' & x"47";
  tmp(325) := 				STA & "00" & '0' & x"20";
  tmp(326) := 				JMP & "00" & '1' & x"48";
  tmp(327) := 					STA & "00" & '0' & x"00";
  tmp(328) := 		STA & "00" & '1' & x"FF";
  tmp(329) := 		LDI & "00" & '0' & x"E0";
  tmp(330) := 		STA & "00" & '1' & x"00";
  tmp(331) := 			LDA & "00" & '1' & x"40";
  tmp(332) := 			LDI & "01" & '0' & x"06";
  tmp(333) := 			CLT & "01" & '1' & x"40";
  tmp(334) := 			JLT & "00" & '1' & x"50";
  tmp(335) := 			JMP & "00" & '1' & x"51";
  tmp(336) := 				LDI & "00" & '0' & x"05";
  tmp(337) := 				STA & "00" & '1' & x"21";
  tmp(338) := 				LDA & "01" & '1' & x"60";
  tmp(339) := 				CEQ & "01" & '0' & x"0A";
  tmp(340) := 				JEQ & "00" & '1' & x"4B";
  tmp(341) := 				STA & "00" & '1' & x"FF";
  tmp(342) := 				LDA & "01" & '0' & x"17";
  tmp(343) := 				CEQ & "01" & '0' & x"0B";
  tmp(344) := 				JEQ & "00" & '1' & x"5B";
  tmp(345) := 				STA & "00" & '0' & x"1F";
  tmp(346) := 				JMP & "00" & '1' & x"5D";
  tmp(347) := 					STA & "00" & '0' & x"32";
  tmp(348) := 					LDA & "11" & '0' & x"32";
  tmp(349) := 		STA & "00" & '1' & x"FF";
  tmp(350) := 		LDI & "00" & '0' & x"F0";
  tmp(351) := 		STA & "00" & '1' & x"00";
  tmp(352) := 			LDA & "00" & '1' & x"40";
  tmp(353) := 			LDI & "01" & '0' & x"0A";
  tmp(354) := 			CLT & "01" & '1' & x"40";
  tmp(355) := 			JLT & "00" & '1' & x"65";
  tmp(356) := 			JMP & "00" & '1' & x"66";
  tmp(357) := 				LDI & "00" & '0' & x"09";
  tmp(358) := 				STA & "00" & '1' & x"20";
  tmp(359) := 				LDA & "01" & '1' & x"60";
  tmp(360) := 				CEQ & "01" & '0' & x"0A";
  tmp(361) := 				JEQ & "00" & '1' & x"60";
  tmp(362) := 				STA & "00" & '1' & x"FF";
  tmp(363) := 				LDA & "01" & '0' & x"17";
  tmp(364) := 				CEQ & "01" & '0' & x"0B";
  tmp(365) := 				JEQ & "00" & '1' & x"70";
  tmp(366) := 				STA & "00" & '0' & x"1E";
  tmp(367) := 				JMP & "00" & '1' & x"72";
  tmp(368) := 					STA & "00" & '0' & x"32";
  tmp(369) := 					LDA & "10" & '0' & x"32";
  tmp(370) := 				LDI & "00" & '0' & x"00";
  tmp(371) := 				LDI & "01" & '0' & x"00";
  tmp(372) := 				STA & "00" & '1' & x"00";
  tmp(373) := 				STA & "00" & '1' & x"01";
  tmp(374) := 				STA & "00" & '1' & x"02";
  tmp(375) := 				RET & "00" & '0' & x"00";
  tmp(376) := 	STA & "00" & '1' & x"FD";
  tmp(377) := 	LDI & "10" & '0' & x"00";
  tmp(378) := 	STA & "10" & '0' & x"00";
  tmp(379) := 	STA & "10" & '0' & x"01";
  tmp(380) := 	STA & "10" & '0' & x"02";
  tmp(381) := 	STA & "10" & '0' & x"03";
  tmp(382) := 	LDI & "11" & '0' & x"01";
  tmp(383) := 	STA & "11" & '0' & x"14";
  tmp(384) := 	LDI & "11" & '0' & x"00";
  tmp(385) := 	RET & "00" & '0' & x"00";
  tmp(386) := 	STA & "00" & '1' & x"FC";
  tmp(387) := 	LDA & "01" & '0' & x"14";
  tmp(388) := 	CEQ & "01" & '0' & x"0B";
  tmp(389) := 	JEQ & "00" & '1' & x"87";
  tmp(390) := 	RET & "00" & '0' & x"00";
  tmp(391) := 		SOMA & "10" & '0' & x"0B";
  tmp(392) := 		CEQ & "10" & '0' & x"0C";
  tmp(393) := 		JEQ & "00" & '1' & x"8B";
  tmp(394) := 		RET & "00" & '0' & x"00";
  tmp(395) := 			SOMA & "11" & '0' & x"0B";
  tmp(396) := 			CEQ & "11" & '0' & x"0D";
  tmp(397) := 			LDI & "10" & '0' & x"00";
  tmp(398) := 			JEQ & "00" & '1' & x"90";
  tmp(399) := 			RET & "00" & '0' & x"00";
  tmp(400) := 				LDI & "00" & '0' & x"01";
  tmp(401) := 				SOMA & "00" & '0' & x"00";
  tmp(402) := 				LDI & "11" & '0' & x"00";
  tmp(403) := 				CEQ & "00" & '0' & x"0C";
  tmp(404) := 				JEQ & "00" & '1' & x"97";
  tmp(405) := 				STA & "00" & '0' & x"00";
  tmp(406) := 				RET & "00" & '0' & x"00";
  tmp(407) := 					LDI & "00" & '0' & x"00";
  tmp(408) := 					STA & "00" & '0' & x"00";
  tmp(409) := 					LDI & "00" & '0' & x"01";
  tmp(410) := 					SOMA & "00" & '0' & x"01";
  tmp(411) := 					CEQ & "00" & '0' & x"0D";
  tmp(412) := 					JEQ & "00" & '1' & x"9F";
  tmp(413) := 					STA & "00" & '0' & x"01";
  tmp(414) := 					RET & "00" & '0' & x"00";
  tmp(415) := 						LDI & "00" & '0' & x"00";
  tmp(416) := 						STA & "00" & '0' & x"01";
  tmp(417) := 						LDI & "00" & '0' & x"01";
  tmp(418) := 						SOMA & "00" & '0' & x"02";
  tmp(419) := 						CEQ & "00" & '0' & x"0C";
  tmp(420) := 						JEQ & "00" & '1' & x"A7";
  tmp(421) := 						STA & "00" & '0' & x"02";
  tmp(422) := 						JMP & "00" & '1' & x"AC";
  tmp(423) := 							LDI & "00" & '0' & x"00";
  tmp(424) := 							STA & "00" & '0' & x"02";
  tmp(425) := 							LDI & "00" & '0' & x"01";
  tmp(426) := 							SOMA & "00" & '0' & x"03";
  tmp(427) := 							STA & "00" & '0' & x"03";
  tmp(428) := 			LDA & "00" & '0' & x"15";
  tmp(429) := 			CEQ & "00" & '0' & x"0A";
  tmp(430) := 			JEQ & "00" & '1' & x"BB";
  tmp(431) := 			LDA & "00" & '0' & x"02";
  tmp(432) := 			CEQ & "00" & '0' & x"0E";
  tmp(433) := 			JEQ & "00" & '1' & x"B3";
  tmp(434) := 			RET & "00" & '0' & x"00";
  tmp(435) := 					LDA & "00" & '0' & x"03";
  tmp(436) := 					CEQ & "00" & '0' & x"0F";
  tmp(437) := 					JEQ & "00" & '1' & x"B7";
  tmp(438) := 					RET & "00" & '0' & x"00";
  tmp(439) := 							LDI & "00" & '0' & x"00";
  tmp(440) := 							STA & "00" & '0' & x"02";
  tmp(441) := 							STA & "00" & '0' & x"03";
  tmp(442) := 							RET & "00" & '0' & x"00";
  tmp(443) := 				LDA & "00" & '0' & x"02";
  tmp(444) := 				CEQ & "00" & '0' & x"0F";
  tmp(445) := 				JEQ & "00" & '1' & x"BF";
  tmp(446) := 				RET & "00" & '0' & x"00";
  tmp(447) := 						LDA & "00" & '0' & x"03";
  tmp(448) := 						CEQ & "00" & '0' & x"0B";
  tmp(449) := 						JEQ & "00" & '1' & x"C3";
  tmp(450) := 						RET & "00" & '0' & x"00";
  tmp(451) := 								LDI & "00" & '0' & x"00";
  tmp(452) := 								STA & "00" & '0' & x"02";
  tmp(453) := 								STA & "00" & '0' & x"03";
  tmp(454) := 								LDA & "00" & '0' & x"16";
  tmp(455) := 								CEQ & "00" & '0' & x"0A";
  tmp(456) := 								JEQ & "00" & '1' & x"CC";
  tmp(457) := 								LDI & "00" & '0' & x"00";
  tmp(458) := 								STA & "00" & '0' & x"16";
  tmp(459) := 								RET & "00" & '0' & x"00";
  tmp(460) := 										LDI & "00" & '0' & x"01";
  tmp(461) := 										STA & "00" & '0' & x"16";
  tmp(462) := 										RET & "00" & '0' & x"00";
  tmp(463) := 	STA & "10" & '1' & x"20";
  tmp(464) := 	STA & "11" & '1' & x"21";
  tmp(465) := 	LDA & "01" & '0' & x"00";
  tmp(466) := 	STA & "01" & '1' & x"22";
  tmp(467) := 	LDA & "01" & '0' & x"01";
  tmp(468) := 	STA & "01" & '1' & x"23";
  tmp(469) := 	LDA & "01" & '0' & x"02";
  tmp(470) := 	STA & "01" & '1' & x"24";
  tmp(471) := 	LDA & "01" & '0' & x"03";
  tmp(472) := 	STA & "01" & '1' & x"25";
  tmp(473) := 	LDA & "01" & '0' & x"15";
  tmp(474) := 	STA & "01" & '1' & x"00";
  tmp(475) := 	LDA & "01" & '0' & x"16";
  tmp(476) := 	STA & "01" & '1' & x"02";
  tmp(477) := 	RET & "00" & '0' & x"00";
  tmp(478) := 	CEQ & "10" & '0' & x"1E";
  tmp(479) := 	JEQ & "00" & '1' & x"E1";
  tmp(480) := 	RET & "00" & '0' & x"00";
  tmp(481) := 		CEQ & "11" & '0' & x"1F";
  tmp(482) := 		JEQ & "00" & '1' & x"E4";
  tmp(483) := 		RET & "00" & '0' & x"00";
  tmp(484) := 			LDA & "00" & '0' & x"00";
  tmp(485) := 			CEQ & "00" & '0' & x"20";
  tmp(486) := 			JEQ & "00" & '1' & x"E8";
  tmp(487) := 			RET & "00" & '0' & x"00";
  tmp(488) := 				LDA & "00" & '0' & x"01";
  tmp(489) := 				CEQ & "00" & '0' & x"21";
  tmp(490) := 				JEQ & "00" & '1' & x"EC";
  tmp(491) := 				RET & "00" & '0' & x"00";
  tmp(492) := 					LDA & "00" & '0' & x"02";
  tmp(493) := 					CEQ & "00" & '0' & x"22";
  tmp(494) := 					JEQ & "00" & '1' & x"F0";
  tmp(495) := 					RET & "00" & '0' & x"00";
  tmp(496) := 						LDA & "00" & '0' & x"03";
  tmp(497) := 						CEQ & "00" & '0' & x"23";
  tmp(498) := 						JEQ & "00" & '1' & x"F4";
  tmp(499) := 						RET & "00" & '0' & x"00";
  tmp(500) := 							LDI & "00" & '0' & x"01";
  tmp(501) := 							STA & "00" & '1' & x"01";
  tmp(502) := 							LDI & "00" & '0' & x"00";
  tmp(503) := 							RET & "00" & '0' & x"00";
        
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;